/*
 * Copyright (c) 2024 Renaldas Zioma
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module atari2600 (
  input wire          clk,
  input wire          reset,
  input wire          system_enable,
  
  input wire   [3:0]  input_switches,
  input wire   [6:0]  input_joystick_0,
  input wire   [6:0]  input_joystick_1,
  input wire   [7:0]  input_paddle_0,
  input wire   [7:0]  input_paddle_1,
  input wire   [7:0]  input_paddle_2,
  input wire   [7:0]  input_paddle_3,

  output wire         rom_read,
  output wire         rom_cycle, // @TODO: this needs to be rethought or atleast better named
  output wire [11:0]  rom_address,
  input  wire  [7:0]  rom_data,
  
  output wire  [6:0]  video,
  output wire  [7:0]  xpos,
  output wire  [8:0]  ypos,
  output wire         vsync,
  output wire         vblank,
  output wire         vwrite,

  output wire  [4:0]  audio
);
  wire _unused_ok = &{input_joystick_1, input_paddle_0, input_paddle_1, input_paddle_2, input_paddle_3};

  assign video = tia_video_out;
  assign audio = tia_audio_l + tia_audio_r;
  
  // Atari 2600 Clocks
  // Video Color Clock: 3.579545 MHz (NTSC), 3.546894 MHz (PAL)
  // CPU Machine Clock: 1.193182 MHz (NTSC), 1.182298 MHz (PAL)
  // The CPU Clock is derived from Video clock divided by three.
  // One color clock = 1 pixel. One machine clock = 3 pixels.
  // pixel ~1:7  VGA clock
  // CPU   ~1:21 VGA clock

  // ===============================================================
  // TIA/PIA/CPU enable strobes/signal generation
  // ===============================================================

  reg  [8:0] clk_counter;
  always @(posedge clk) begin
    if (reset)
      clk_counter <= 0;
    else if (system_enable) begin
      if (clk_counter >= 3)
        clk_counter <= 0;
      else
        clk_counter <= clk_counter + 1;
    end
  end

  // Strobes (enable) signals emulate the 3 clocks of the Atari 2600 system:
  // tia_enable - XTAL 3.57 MHz system master clock / NTSC clock
  // cpu_enable - PHI0 generated by TIA and driving CPU clock
  // pia_enable - PHI2 generated by CPU and driving PIA clock
  wire tia_enable = system_enable && (clk_counter == 0 || 
                                      clk_counter == 2 ||
                                      clk_counter == 3);
  wire cpu_enable = system_enable &&  clk_counter == 1; // TIA & CPU must tick on a different cycle, otherwise player sprites jitter
  wire pia_enable = system_enable &&  clk_counter == 2;

  assign rom_cycle = (clk_counter == 1);

  // ===============================================================
  // TIA/PIA/RAM/CPU chips
  // ===============================================================
  wire [15:0] address_bus_w;
  reg  [15:0] address_bus_r;
  wire [15:0] address_bus = cpu_enable ? address_bus_w : address_bus_r;
  reg  [7:0] data_in; // register - because that's how Arlet Otten's 6502 impl wants it
  wire [7:0] data_out;
  wire write_enable;
  reg stall_cpu;

  always @(posedge clk)
    if (reset)
      address_bus_r <= 0;
    else
      address_bus_r <= address_bus;

  cpu cpu(
    .clk(clk),
    .reset(reset),
    .AB(address_bus_w),
    .DI(data_in),
    .DO(data_out),
    .WE(write_enable),
    .IRQ(1'b0),  // pins are not inverted in Arlet Otten's 6502 impl
    .NMI(1'b0),  // pins are not inverted in Arlet Otten's 6502 impl
    .RDY(cpu_enable && !stall_cpu)
    );

  wire [3:0] tia_audio_l;
  wire [3:0] tia_audio_r;
  wire [7:0] tia_data_in = data_out;
  reg  [7:0] tia_data_out;
  reg  [6:0] tia_video_out;
  wire [8:0] tia_ypos;  // used to syncronize VGA & TIA frames

  tia tia (
    .clk_i(clk),
    .rst_i(reset),
    .stb_i(tia_cs && cpu_enable),
    .we_i(write_enable),
    .adr_i(address_bus[5:0]),
    .dat_i(tia_data_in),
    .dat_o(tia_data_out),
    .buttons(input_joystick_0),
    .pot(input_paddle_0),
    .audio_left(tia_audio_l),
    .audio_right(tia_audio_r),
    .stall_cpu(stall_cpu),
    .enable_i(tia_enable),
    .cpu_enable_i(cpu_enable),
    .vid_out(tia_video_out),
    .vid_xpos(xpos),
    .vid_ypos(ypos),
    .vid_vblank(vblank),
    .vid_vsync(vsync),
    .vid_wr(video_write),
    .pal(1'b0)  // currently only NSTC is supported
  );

  wire [7:0] pia_data_in = data_out;
  reg  [7:0] pia_data_out;

  pia pia (
    .clk_i(clk),
    .rst_i(reset),
    .enable_i(pia_enable),
    .stb_i(pia_cs && cpu_enable),
    .we_i(write_enable),
    .adr_i(address_bus[6:0]),
    .dat_i(pia_data_in),
    .dat_o(pia_data_out),
    .buttons(input_joystick_0),
    .sw(input_switches)
  );

  reg [7:0] ram [ 127:0]; // Built-in RAM (part of PIA/RIOT chip): 128 bytes
  reg [7:0] ram_data;     // registering this makes yosys iCE40 BRAM inference happy

  // ===============================================================
  // Memory Map
  // ===============================================================

  // All memory is mirrored in steps of 2000h
  // TIA Write Mirrors (Step 40h,100h)
  // TIA Read Mirrors (Step 10h,100h)
  // PIA I/O Mirrors (Step 2h,8h,100h,400h)
  // PIA RAM Mirrors (Step 100h,400h)
  // 0000-002C  TIA Write
  // 0000-000D  TIA Read
  // 0080-00FF  PIA RAM (128 bytes)
  // 0280-0297  PIA Reads & Writes
  // F000-FFFF  Cartridge Memory (4 Kbytes area)

  // From Atari 2600 schematics:
  // - TIA select = ~A12 (-> TIA /CS0) & ~A7 (-> TIA /CS3)
  // - PIA select = ~A12 (-> PIA /CS2) &  A7 (-> PIA  CS1) &  A9 ('1' -> PIA RS)
  // - RAM select = ~A12 (-> PIA /CS2) &  A7 (-> PIA  CS1) & ~A9 ('0' -> PIA RS)

  wire rom_cs = (address_bus[12] == 1);
  wire tia_cs = (address_bus[12] == 0 && address_bus[7] == 0);
  wire pia_cs = (address_bus[12] == 0 && address_bus[7] == 1 && address_bus[9] == 1);
  wire ram_cs = (address_bus[12] == 0 && address_bus[7] == 1 && address_bus[9] == 0);

  assign rom_read = cpu_enable && !stall_cpu && rom_cs;
  assign rom_address = address_bus[11:0];

  always @(posedge clk) begin
    // CPU writes
    if (cpu_enable && write_enable && ram_cs) ram[address_bus[6:0]] <= data_out;
    // if (~write_enable && ram_cs)              ram_data <= ram[address_bus[6:0]]; 

    // CPU reads
    if (~write_enable &&
        ram_cs) data_in <= ram[address_bus[6:0]];
    if (rom_cs) data_in <= rom_data;
    if (tia_cs) data_in <= tia_data_out;
    if (pia_cs) data_in <= pia_data_out;
  end

endmodule
