`ifndef HVSYNC_GENERATOR_H
`define HVSYNC_GENERATOR_H

/*
Video sync generator, used to drive a VGA monitor.
Timing from: https://en.wikipedia.org/wiki/Video_Graphics_Array
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
*/

module vga_640x480_25MHz_hvsync_generator(
  input clk,
  input reset,
  output reg hsync,
  output reg vsync,
  output display_on,
  output reg [9:0] hpos,
  output reg [9:0] vpos
);
  vga_hvsync_generator vga (
    .clk, .reset, .hsync, .vsync, .display_on, .hpos, .vpos
  );
endmodule

module vga_640x480_50MHz_hvsync_generator(
  input clk,
  input reset,
  output reg hsync,
  output reg vsync,
  output display_on,
  output reg [9:0] hpos,
  output reg [9:0] vpos
);
  reg sub_pixel;
  vga_hvsync_generator #(
    .H_DISPLAY(640 * 2),  // horizontal display width
    .H_BACK   ( 48 * 2),  // horizontal left border (back porch)
    .H_FRONT  ( 16 * 2),  // horizontal right border (front porch)
    .H_SYNC   ( 96 * 2)   // horizontal sync width
  ) vga (
    .clk, .reset, .hsync, .vsync, .display_on, .vpos,
    .hpos      ({hpos, sub_pixel})
  );
endmodule

module vga_1280x480_50MHz_hvsync_generator(
  input clk,
  input reset,
  output reg hsync,
  output reg vsync,
  output display_on,
  output reg [10:0] hpos,
  output reg [ 9:0] vpos
);
  vga_hvsync_generator #(
    .H_DISPLAY(640 * 2),  // horizontal display width
    .H_BACK   ( 48 * 2),  // horizontal left border (back porch)
    .H_FRONT  ( 16 * 2),  // horizontal right border (front porch)
    .H_SYNC   ( 96 * 2)   // horizontal sync width
  ) vga (
    .clk, .reset, .hsync, .vsync, .display_on, .hpos, .vpos
  );
endmodule

module vga_hvsync_generator #(
  // declarations for TV-simulator sync parameters
  // horizontal constants
  parameter H_DISPLAY       = 640, // horizontal display width
  parameter H_BACK          =  48, // horizontal left border (back porch)
  parameter H_FRONT         =  16, // horizontal right border (front porch)
  parameter H_SYNC          =  96, // horizontal sync width
  // vertical constants
  parameter V_DISPLAY       = 480, // vertical display height
  parameter V_TOP           =  33, // vertical top border
  parameter V_BOTTOM        =  10, // vertical bottom border
  parameter V_SYNC          =   2  // vertical sync # lines
) ( clk, reset, hsync, vsync, display_on, hpos, vpos);

  input clk;
  input reset;
  output reg hsync, vsync;
  output display_on;
  output reg [$clog2(H_MAX)-1:0] hpos;
  output reg [$clog2(V_MAX)-1:0] vpos;

  // derived constants
  parameter H_SYNC_START    = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END      = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX           = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START    = 0;
  parameter V_SYNC_END      = 0 + V_SYNC - 1;
  parameter V_MAX           = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

  wire hmaxxed = (hpos == H_MAX) || reset;  // set when hpos is maximum
  wire vmaxxed = (vpos == V_MAX) || reset;  // set when vpos is maximum
  
  // horizontal position counter
  always @(posedge clk)
  begin
    hsync <= (hpos>=H_SYNC_START && hpos<=H_SYNC_END);
    if (hmaxxed)
      hpos <= 0;
    else
      hpos <= hpos + 1;
  end

  // vertical position counter
  always @(posedge clk)
  begin
    vsync <= (                      vpos<=V_SYNC_END);
    if (hmaxxed)
      if (vmaxxed)
        vpos <= 0;
      else
        vpos <= vpos + 1;
  end
  
  // display_on is set when beam is in "safe" visible frame
  assign display_on = (hpos<H_DISPLAY) && (vpos<V_DISPLAY);

endmodule

`endif
